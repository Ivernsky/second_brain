module TOP;
  wire [1:0] w1;
  wire w2, w3;
  wire w4[7:0][255:0];
  wire ws[3:0];
endmodule


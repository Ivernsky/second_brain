
module top;
  bind top.k0 m i0();
  k k0();
endmodule

module m;
endmodule

module k;
endmodule

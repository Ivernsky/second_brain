module top;
  m #(2) i0();
endmodule

module m();
  parameter P = 1;
endmodule 

module MOD;
  wire a;
endmodule

module test (a, b, c);
  input a, b;
  output c;
 
  and and_gate (c, a, b);
endmodule

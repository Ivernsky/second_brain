module top;
  dly u_dlu();
  FD1 u_fd1();
endmodule

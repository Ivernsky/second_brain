module test (a, b, c);
/* line 2 will be replaced */
  input a, b;
  output c;
  wire c;
 
  and and_gate (c, a, b);
endmodule

module top;
  wire [3:0] a = 4'b1110; // 3-bit net with identifier "a"
  wire \b[3:0]  = 1'b1;    // 1-bit net with escape identifier "\b[3:0] "
endmodule

module top;
  logic a;
  reg c;
endmodule

module myand (a, b, c);
  input a, b;
  output c;
  wire c;
 
  and myandgate (c, a, b);
endmodule

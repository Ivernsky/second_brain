module TOP;
endmodule


module top;
  parameter pi = 3.14;
endmodule

module top;
  wire [0:3] a, b;
  wire c;
  assign b = a;
  assign c = a[0];
endmodule 

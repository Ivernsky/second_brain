module TOP;
  logic a, b, c;
  
  always@(posedge a) begin
    b<=c;
  end 
endmodule


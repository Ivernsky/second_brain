module top;
  typedef logic T1;
endmodule

module top;
  wire a, b;
  assign a = b;
endmodule

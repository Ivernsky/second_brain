module TOP;
  wire a, b;

  MOD i0( a, b );
endmodule

module MOD( input a, b );
endmodule

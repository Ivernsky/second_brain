module MOD;
endmodule

module TOP;
  MOD inst();
  MOD inst2 [3:0] ();
endmodule



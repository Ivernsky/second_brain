module test (a, b, c);
  input a, b;;
  output c;
  wire c;
 
  and and_gate (c, a, b);
endmodule

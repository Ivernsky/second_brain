module MOD;
  wire a, b;
  assign a = b;
endmodule


module MOD;
  logic a, b;
endmodule

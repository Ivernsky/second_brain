module top;
  dly u_dly();
  FD1 u_fd1();
endmodule

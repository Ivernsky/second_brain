package pkg;
  bit a;
endpackage

module TOP;
endmodule


module test;
parameter PARAM_BIN     = 5'bxxz10;
parameter PARAM_DEC     = 10'd123;
parameter PARAM_OCT     = 24'o7777_7777;
parameter PARAM_HEX     = 32'hffff_ffff;
parameter PARAM_INTEGER = 111004;
parameter PARAM_REAL    = 1.25;
parameter PARAM_STRING  = "springsoft";
parameter PARAM_UNBOUND = 'x;
endmodule

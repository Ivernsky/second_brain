module TOP;
  MOD i0();
endmodule

module MOD;
endmodule


module mem;
endmodule

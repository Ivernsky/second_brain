module MOD;
  wire a;
  logic b;
endmodule

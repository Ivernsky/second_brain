module top;
  cpu i_cpu();
endmodule

module TOP;
  wire a, b;
  assign a = b;
endmodule


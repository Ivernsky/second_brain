module TOP;
  wire ndm_net;
  MOD i0();
endmodule

module MOD;
endmodule


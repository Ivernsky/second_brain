module top;
  wire signed [3:0] a, b, c, d, e, f;
  assign a = b | c;
  assign d = e + f;
endmodule

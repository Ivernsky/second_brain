module top;
  parameter P1 = 1;
  parameter P2 = 2;
endmodule

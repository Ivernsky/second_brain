module TOP;
  MOD #( .P( 2 ), .PT( bit ) ) i0();
endmodule

module MOD;
  parameter P = 1 ;
  parameter type PT = logic;
endmodule


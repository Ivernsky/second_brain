module TOP;
  wire [4:0] w1 [2:0];
endmodule

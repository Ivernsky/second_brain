module TOP;
  logic a, b, c;
  assign a = b ? 1'bz : c;  
endmodule


interface Itf;
endinterface

module TOP;
  Itf i0();
endmodule


module top;
 
parameter P1 = 31;
parameter P2 = 4'b1111;
integer a = P1 - P2 + 3.2 / 2 + P1;

endmodule

module TOP;
  wire a, b;
  MOD ndm_instance( a, b );
endmodule

module MOD( a, b );
  input  a;
  output b;
endmodule


module MOD;
  wor w1 [3:0];
  supply1 sp1;
  wire [2:0] w2 [4:0];
endmodule

module TOP;
  MOD inst();
endmodule

module top;

wire [3:0] w;
wire [1:0] a, b;
assign w = {a, b};

endmodule

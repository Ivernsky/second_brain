module MOD;
  parameter type PT = logic;
endmodule

module TOP;
  parameter P1 = 1;
  MOD i0();
endmodule

module MOD;
  parameter P2 = 2;
endmodule

module TOP;
  parameter P1 = 1;
  MOD i0();
endmodule


module datapath;
endmodule

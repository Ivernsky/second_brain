module top;
  wire [31:0] a, b, c;
  AN2 u1(a,b,c);
endmodule

module top;
  wire a, b, c;
  assign a = b;
  assign b = c;
endmodule

module top;
 
    parameter PARAM_INTEGER = -111004;
    parameter PARAM_BIN = 5'bxxz10;
    parameter PARAM_HEX = 32'hffff_ffff;
    parameter PARAM_OCT = 'o7777_7777_7777;
    parameter PARAM_DEC = 10'sd1023;
    parameter PARAM_REAL = 1.25;
    parameter PARAM_STRING = "springsoft";
 
endmodule

module TOP;
  wire a, b;
  MOD ndm_instance( a, b );
endmodule

module MOD( input a, b );
endmodule


module top;
  wire a;
  m i0( a );
endmodule

module m( input a );
endmodule 


module top;
  wire  w1, w2, w3;
  assign w1 = w2 & w3;
endmodule

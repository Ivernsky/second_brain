module mm;
   reg mr;
endmodule
 
module top;
    bit [3:0] r;
    mm mArr [1:0] ();
endmodule

module cpu;
  alu i1();
  mem i2();
  datapath i3();
endmodule

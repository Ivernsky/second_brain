module top;
    bit [5:0] r;
endmodule

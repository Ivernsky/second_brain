module MOD;
  logic a;
endmodule
